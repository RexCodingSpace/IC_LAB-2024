# 
#              Synchronous High Speed Single Port SRAM Compiler 
# 
#                    UMC 0.18um GenericII Logic Process
#    __________________________________________________________________________
# 
# 
#      (C) Copyright 2002-2009 Faraday Technology Corp. All Rights Reserved.
#    
#    This source code is an unpublished work belongs to Faraday Technology
#    Corp.  It is considered a trade secret and is not to be divulged or
#    used by parties who have not received written authorization from
#    Faraday Technology Corp.
#    
#    Faraday's home page can be found at:
#    http://www.faraday-tech.com/
#   
#       Module Name      : MEM1_1
#       Words            : 512
#       Bits             : 16
#       Byte-Write       : 1
#       Aspect Ratio     : 1
#       Output Loading   : 0.05  (pf)
#       Data Slew        : 0.02  (ns)
#       CK Slew          : 0.02  (ns)
#       Power Ring Width : 2  (um)
# 
# -----------------------------------------------------------------------------
# 
#       Library          : FSA0M_A
#       Memaker          : 200901.2.1
#       Date             : 2024/10/10 15:39:33
# 
# -----------------------------------------------------------------------------


NAMESCASESENSITIVE ON ;
MACRO MEM1_1
CLASS BLOCK ;
FOREIGN MEM1_1 0.000 0.000 ;
ORIGIN 0.000 0.000 ;
SIZE 326.740 BY 294.000 ;
SYMMETRY x y r90 ;
SITE core ;
PIN VCC
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
 PORT
  LAYER ME4 ;
  RECT 325.620 282.580 326.740 285.820 ;
  LAYER ME3 ;
  RECT 325.620 282.580 326.740 285.820 ;
  LAYER ME2 ;
  RECT 325.620 282.580 326.740 285.820 ;
  LAYER ME1 ;
  RECT 325.620 282.580 326.740 285.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.620 274.740 326.740 277.980 ;
  LAYER ME3 ;
  RECT 325.620 274.740 326.740 277.980 ;
  LAYER ME2 ;
  RECT 325.620 274.740 326.740 277.980 ;
  LAYER ME1 ;
  RECT 325.620 274.740 326.740 277.980 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.620 266.900 326.740 270.140 ;
  LAYER ME3 ;
  RECT 325.620 266.900 326.740 270.140 ;
  LAYER ME2 ;
  RECT 325.620 266.900 326.740 270.140 ;
  LAYER ME1 ;
  RECT 325.620 266.900 326.740 270.140 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.620 259.060 326.740 262.300 ;
  LAYER ME3 ;
  RECT 325.620 259.060 326.740 262.300 ;
  LAYER ME2 ;
  RECT 325.620 259.060 326.740 262.300 ;
  LAYER ME1 ;
  RECT 325.620 259.060 326.740 262.300 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.620 251.220 326.740 254.460 ;
  LAYER ME3 ;
  RECT 325.620 251.220 326.740 254.460 ;
  LAYER ME2 ;
  RECT 325.620 251.220 326.740 254.460 ;
  LAYER ME1 ;
  RECT 325.620 251.220 326.740 254.460 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.620 243.380 326.740 246.620 ;
  LAYER ME3 ;
  RECT 325.620 243.380 326.740 246.620 ;
  LAYER ME2 ;
  RECT 325.620 243.380 326.740 246.620 ;
  LAYER ME1 ;
  RECT 325.620 243.380 326.740 246.620 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.620 204.180 326.740 207.420 ;
  LAYER ME3 ;
  RECT 325.620 204.180 326.740 207.420 ;
  LAYER ME2 ;
  RECT 325.620 204.180 326.740 207.420 ;
  LAYER ME1 ;
  RECT 325.620 204.180 326.740 207.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.620 196.340 326.740 199.580 ;
  LAYER ME3 ;
  RECT 325.620 196.340 326.740 199.580 ;
  LAYER ME2 ;
  RECT 325.620 196.340 326.740 199.580 ;
  LAYER ME1 ;
  RECT 325.620 196.340 326.740 199.580 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.620 188.500 326.740 191.740 ;
  LAYER ME3 ;
  RECT 325.620 188.500 326.740 191.740 ;
  LAYER ME2 ;
  RECT 325.620 188.500 326.740 191.740 ;
  LAYER ME1 ;
  RECT 325.620 188.500 326.740 191.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.620 180.660 326.740 183.900 ;
  LAYER ME3 ;
  RECT 325.620 180.660 326.740 183.900 ;
  LAYER ME2 ;
  RECT 325.620 180.660 326.740 183.900 ;
  LAYER ME1 ;
  RECT 325.620 180.660 326.740 183.900 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.620 172.820 326.740 176.060 ;
  LAYER ME3 ;
  RECT 325.620 172.820 326.740 176.060 ;
  LAYER ME2 ;
  RECT 325.620 172.820 326.740 176.060 ;
  LAYER ME1 ;
  RECT 325.620 172.820 326.740 176.060 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.620 164.980 326.740 168.220 ;
  LAYER ME3 ;
  RECT 325.620 164.980 326.740 168.220 ;
  LAYER ME2 ;
  RECT 325.620 164.980 326.740 168.220 ;
  LAYER ME1 ;
  RECT 325.620 164.980 326.740 168.220 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.620 125.780 326.740 129.020 ;
  LAYER ME3 ;
  RECT 325.620 125.780 326.740 129.020 ;
  LAYER ME2 ;
  RECT 325.620 125.780 326.740 129.020 ;
  LAYER ME1 ;
  RECT 325.620 125.780 326.740 129.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.620 117.940 326.740 121.180 ;
  LAYER ME3 ;
  RECT 325.620 117.940 326.740 121.180 ;
  LAYER ME2 ;
  RECT 325.620 117.940 326.740 121.180 ;
  LAYER ME1 ;
  RECT 325.620 117.940 326.740 121.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.620 110.100 326.740 113.340 ;
  LAYER ME3 ;
  RECT 325.620 110.100 326.740 113.340 ;
  LAYER ME2 ;
  RECT 325.620 110.100 326.740 113.340 ;
  LAYER ME1 ;
  RECT 325.620 110.100 326.740 113.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.620 102.260 326.740 105.500 ;
  LAYER ME3 ;
  RECT 325.620 102.260 326.740 105.500 ;
  LAYER ME2 ;
  RECT 325.620 102.260 326.740 105.500 ;
  LAYER ME1 ;
  RECT 325.620 102.260 326.740 105.500 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.620 94.420 326.740 97.660 ;
  LAYER ME3 ;
  RECT 325.620 94.420 326.740 97.660 ;
  LAYER ME2 ;
  RECT 325.620 94.420 326.740 97.660 ;
  LAYER ME1 ;
  RECT 325.620 94.420 326.740 97.660 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.620 86.580 326.740 89.820 ;
  LAYER ME3 ;
  RECT 325.620 86.580 326.740 89.820 ;
  LAYER ME2 ;
  RECT 325.620 86.580 326.740 89.820 ;
  LAYER ME1 ;
  RECT 325.620 86.580 326.740 89.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.620 47.380 326.740 50.620 ;
  LAYER ME3 ;
  RECT 325.620 47.380 326.740 50.620 ;
  LAYER ME2 ;
  RECT 325.620 47.380 326.740 50.620 ;
  LAYER ME1 ;
  RECT 325.620 47.380 326.740 50.620 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.620 39.540 326.740 42.780 ;
  LAYER ME3 ;
  RECT 325.620 39.540 326.740 42.780 ;
  LAYER ME2 ;
  RECT 325.620 39.540 326.740 42.780 ;
  LAYER ME1 ;
  RECT 325.620 39.540 326.740 42.780 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.620 31.700 326.740 34.940 ;
  LAYER ME3 ;
  RECT 325.620 31.700 326.740 34.940 ;
  LAYER ME2 ;
  RECT 325.620 31.700 326.740 34.940 ;
  LAYER ME1 ;
  RECT 325.620 31.700 326.740 34.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.620 23.860 326.740 27.100 ;
  LAYER ME3 ;
  RECT 325.620 23.860 326.740 27.100 ;
  LAYER ME2 ;
  RECT 325.620 23.860 326.740 27.100 ;
  LAYER ME1 ;
  RECT 325.620 23.860 326.740 27.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.620 16.020 326.740 19.260 ;
  LAYER ME3 ;
  RECT 325.620 16.020 326.740 19.260 ;
  LAYER ME2 ;
  RECT 325.620 16.020 326.740 19.260 ;
  LAYER ME1 ;
  RECT 325.620 16.020 326.740 19.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.620 8.180 326.740 11.420 ;
  LAYER ME3 ;
  RECT 325.620 8.180 326.740 11.420 ;
  LAYER ME2 ;
  RECT 325.620 8.180 326.740 11.420 ;
  LAYER ME1 ;
  RECT 325.620 8.180 326.740 11.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 282.580 1.120 285.820 ;
  LAYER ME3 ;
  RECT 0.000 282.580 1.120 285.820 ;
  LAYER ME2 ;
  RECT 0.000 282.580 1.120 285.820 ;
  LAYER ME1 ;
  RECT 0.000 282.580 1.120 285.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 274.740 1.120 277.980 ;
  LAYER ME3 ;
  RECT 0.000 274.740 1.120 277.980 ;
  LAYER ME2 ;
  RECT 0.000 274.740 1.120 277.980 ;
  LAYER ME1 ;
  RECT 0.000 274.740 1.120 277.980 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 266.900 1.120 270.140 ;
  LAYER ME3 ;
  RECT 0.000 266.900 1.120 270.140 ;
  LAYER ME2 ;
  RECT 0.000 266.900 1.120 270.140 ;
  LAYER ME1 ;
  RECT 0.000 266.900 1.120 270.140 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 259.060 1.120 262.300 ;
  LAYER ME3 ;
  RECT 0.000 259.060 1.120 262.300 ;
  LAYER ME2 ;
  RECT 0.000 259.060 1.120 262.300 ;
  LAYER ME1 ;
  RECT 0.000 259.060 1.120 262.300 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 251.220 1.120 254.460 ;
  LAYER ME3 ;
  RECT 0.000 251.220 1.120 254.460 ;
  LAYER ME2 ;
  RECT 0.000 251.220 1.120 254.460 ;
  LAYER ME1 ;
  RECT 0.000 251.220 1.120 254.460 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 243.380 1.120 246.620 ;
  LAYER ME3 ;
  RECT 0.000 243.380 1.120 246.620 ;
  LAYER ME2 ;
  RECT 0.000 243.380 1.120 246.620 ;
  LAYER ME1 ;
  RECT 0.000 243.380 1.120 246.620 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 204.180 1.120 207.420 ;
  LAYER ME3 ;
  RECT 0.000 204.180 1.120 207.420 ;
  LAYER ME2 ;
  RECT 0.000 204.180 1.120 207.420 ;
  LAYER ME1 ;
  RECT 0.000 204.180 1.120 207.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 196.340 1.120 199.580 ;
  LAYER ME3 ;
  RECT 0.000 196.340 1.120 199.580 ;
  LAYER ME2 ;
  RECT 0.000 196.340 1.120 199.580 ;
  LAYER ME1 ;
  RECT 0.000 196.340 1.120 199.580 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 188.500 1.120 191.740 ;
  LAYER ME3 ;
  RECT 0.000 188.500 1.120 191.740 ;
  LAYER ME2 ;
  RECT 0.000 188.500 1.120 191.740 ;
  LAYER ME1 ;
  RECT 0.000 188.500 1.120 191.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 180.660 1.120 183.900 ;
  LAYER ME3 ;
  RECT 0.000 180.660 1.120 183.900 ;
  LAYER ME2 ;
  RECT 0.000 180.660 1.120 183.900 ;
  LAYER ME1 ;
  RECT 0.000 180.660 1.120 183.900 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 172.820 1.120 176.060 ;
  LAYER ME3 ;
  RECT 0.000 172.820 1.120 176.060 ;
  LAYER ME2 ;
  RECT 0.000 172.820 1.120 176.060 ;
  LAYER ME1 ;
  RECT 0.000 172.820 1.120 176.060 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 164.980 1.120 168.220 ;
  LAYER ME3 ;
  RECT 0.000 164.980 1.120 168.220 ;
  LAYER ME2 ;
  RECT 0.000 164.980 1.120 168.220 ;
  LAYER ME1 ;
  RECT 0.000 164.980 1.120 168.220 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER ME3 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER ME2 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER ME1 ;
  RECT 0.000 125.780 1.120 129.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER ME3 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER ME2 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER ME1 ;
  RECT 0.000 117.940 1.120 121.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER ME3 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER ME2 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER ME1 ;
  RECT 0.000 110.100 1.120 113.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER ME3 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER ME2 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER ME1 ;
  RECT 0.000 102.260 1.120 105.500 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER ME3 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER ME2 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER ME1 ;
  RECT 0.000 94.420 1.120 97.660 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER ME3 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER ME2 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER ME1 ;
  RECT 0.000 86.580 1.120 89.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER ME3 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER ME2 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER ME1 ;
  RECT 0.000 47.380 1.120 50.620 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER ME3 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER ME2 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER ME1 ;
  RECT 0.000 39.540 1.120 42.780 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER ME3 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER ME2 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER ME1 ;
  RECT 0.000 31.700 1.120 34.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER ME3 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER ME2 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER ME1 ;
  RECT 0.000 23.860 1.120 27.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER ME3 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER ME2 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER ME1 ;
  RECT 0.000 16.020 1.120 19.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER ME3 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER ME2 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER ME1 ;
  RECT 0.000 8.180 1.120 11.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 311.640 292.880 315.180 294.000 ;
  LAYER ME3 ;
  RECT 311.640 292.880 315.180 294.000 ;
  LAYER ME2 ;
  RECT 311.640 292.880 315.180 294.000 ;
  LAYER ME1 ;
  RECT 311.640 292.880 315.180 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 302.960 292.880 306.500 294.000 ;
  LAYER ME3 ;
  RECT 302.960 292.880 306.500 294.000 ;
  LAYER ME2 ;
  RECT 302.960 292.880 306.500 294.000 ;
  LAYER ME1 ;
  RECT 302.960 292.880 306.500 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 294.280 292.880 297.820 294.000 ;
  LAYER ME3 ;
  RECT 294.280 292.880 297.820 294.000 ;
  LAYER ME2 ;
  RECT 294.280 292.880 297.820 294.000 ;
  LAYER ME1 ;
  RECT 294.280 292.880 297.820 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 285.600 292.880 289.140 294.000 ;
  LAYER ME3 ;
  RECT 285.600 292.880 289.140 294.000 ;
  LAYER ME2 ;
  RECT 285.600 292.880 289.140 294.000 ;
  LAYER ME1 ;
  RECT 285.600 292.880 289.140 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 276.920 292.880 280.460 294.000 ;
  LAYER ME3 ;
  RECT 276.920 292.880 280.460 294.000 ;
  LAYER ME2 ;
  RECT 276.920 292.880 280.460 294.000 ;
  LAYER ME1 ;
  RECT 276.920 292.880 280.460 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 268.240 292.880 271.780 294.000 ;
  LAYER ME3 ;
  RECT 268.240 292.880 271.780 294.000 ;
  LAYER ME2 ;
  RECT 268.240 292.880 271.780 294.000 ;
  LAYER ME1 ;
  RECT 268.240 292.880 271.780 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 224.840 292.880 228.380 294.000 ;
  LAYER ME3 ;
  RECT 224.840 292.880 228.380 294.000 ;
  LAYER ME2 ;
  RECT 224.840 292.880 228.380 294.000 ;
  LAYER ME1 ;
  RECT 224.840 292.880 228.380 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 216.160 292.880 219.700 294.000 ;
  LAYER ME3 ;
  RECT 216.160 292.880 219.700 294.000 ;
  LAYER ME2 ;
  RECT 216.160 292.880 219.700 294.000 ;
  LAYER ME1 ;
  RECT 216.160 292.880 219.700 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 207.480 292.880 211.020 294.000 ;
  LAYER ME3 ;
  RECT 207.480 292.880 211.020 294.000 ;
  LAYER ME2 ;
  RECT 207.480 292.880 211.020 294.000 ;
  LAYER ME1 ;
  RECT 207.480 292.880 211.020 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 198.800 292.880 202.340 294.000 ;
  LAYER ME3 ;
  RECT 198.800 292.880 202.340 294.000 ;
  LAYER ME2 ;
  RECT 198.800 292.880 202.340 294.000 ;
  LAYER ME1 ;
  RECT 198.800 292.880 202.340 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 190.120 292.880 193.660 294.000 ;
  LAYER ME3 ;
  RECT 190.120 292.880 193.660 294.000 ;
  LAYER ME2 ;
  RECT 190.120 292.880 193.660 294.000 ;
  LAYER ME1 ;
  RECT 190.120 292.880 193.660 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 181.440 292.880 184.980 294.000 ;
  LAYER ME3 ;
  RECT 181.440 292.880 184.980 294.000 ;
  LAYER ME2 ;
  RECT 181.440 292.880 184.980 294.000 ;
  LAYER ME1 ;
  RECT 181.440 292.880 184.980 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 138.040 292.880 141.580 294.000 ;
  LAYER ME3 ;
  RECT 138.040 292.880 141.580 294.000 ;
  LAYER ME2 ;
  RECT 138.040 292.880 141.580 294.000 ;
  LAYER ME1 ;
  RECT 138.040 292.880 141.580 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 129.360 292.880 132.900 294.000 ;
  LAYER ME3 ;
  RECT 129.360 292.880 132.900 294.000 ;
  LAYER ME2 ;
  RECT 129.360 292.880 132.900 294.000 ;
  LAYER ME1 ;
  RECT 129.360 292.880 132.900 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 120.680 292.880 124.220 294.000 ;
  LAYER ME3 ;
  RECT 120.680 292.880 124.220 294.000 ;
  LAYER ME2 ;
  RECT 120.680 292.880 124.220 294.000 ;
  LAYER ME1 ;
  RECT 120.680 292.880 124.220 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 112.000 292.880 115.540 294.000 ;
  LAYER ME3 ;
  RECT 112.000 292.880 115.540 294.000 ;
  LAYER ME2 ;
  RECT 112.000 292.880 115.540 294.000 ;
  LAYER ME1 ;
  RECT 112.000 292.880 115.540 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 103.320 292.880 106.860 294.000 ;
  LAYER ME3 ;
  RECT 103.320 292.880 106.860 294.000 ;
  LAYER ME2 ;
  RECT 103.320 292.880 106.860 294.000 ;
  LAYER ME1 ;
  RECT 103.320 292.880 106.860 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 94.640 292.880 98.180 294.000 ;
  LAYER ME3 ;
  RECT 94.640 292.880 98.180 294.000 ;
  LAYER ME2 ;
  RECT 94.640 292.880 98.180 294.000 ;
  LAYER ME1 ;
  RECT 94.640 292.880 98.180 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 51.240 292.880 54.780 294.000 ;
  LAYER ME3 ;
  RECT 51.240 292.880 54.780 294.000 ;
  LAYER ME2 ;
  RECT 51.240 292.880 54.780 294.000 ;
  LAYER ME1 ;
  RECT 51.240 292.880 54.780 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 42.560 292.880 46.100 294.000 ;
  LAYER ME3 ;
  RECT 42.560 292.880 46.100 294.000 ;
  LAYER ME2 ;
  RECT 42.560 292.880 46.100 294.000 ;
  LAYER ME1 ;
  RECT 42.560 292.880 46.100 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 33.880 292.880 37.420 294.000 ;
  LAYER ME3 ;
  RECT 33.880 292.880 37.420 294.000 ;
  LAYER ME2 ;
  RECT 33.880 292.880 37.420 294.000 ;
  LAYER ME1 ;
  RECT 33.880 292.880 37.420 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 25.200 292.880 28.740 294.000 ;
  LAYER ME3 ;
  RECT 25.200 292.880 28.740 294.000 ;
  LAYER ME2 ;
  RECT 25.200 292.880 28.740 294.000 ;
  LAYER ME1 ;
  RECT 25.200 292.880 28.740 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 16.520 292.880 20.060 294.000 ;
  LAYER ME3 ;
  RECT 16.520 292.880 20.060 294.000 ;
  LAYER ME2 ;
  RECT 16.520 292.880 20.060 294.000 ;
  LAYER ME1 ;
  RECT 16.520 292.880 20.060 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 7.840 292.880 11.380 294.000 ;
  LAYER ME3 ;
  RECT 7.840 292.880 11.380 294.000 ;
  LAYER ME2 ;
  RECT 7.840 292.880 11.380 294.000 ;
  LAYER ME1 ;
  RECT 7.840 292.880 11.380 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 307.300 0.000 310.840 1.120 ;
  LAYER ME3 ;
  RECT 307.300 0.000 310.840 1.120 ;
  LAYER ME2 ;
  RECT 307.300 0.000 310.840 1.120 ;
  LAYER ME1 ;
  RECT 307.300 0.000 310.840 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 285.600 0.000 289.140 1.120 ;
  LAYER ME3 ;
  RECT 285.600 0.000 289.140 1.120 ;
  LAYER ME2 ;
  RECT 285.600 0.000 289.140 1.120 ;
  LAYER ME1 ;
  RECT 285.600 0.000 289.140 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 263.900 0.000 267.440 1.120 ;
  LAYER ME3 ;
  RECT 263.900 0.000 267.440 1.120 ;
  LAYER ME2 ;
  RECT 263.900 0.000 267.440 1.120 ;
  LAYER ME1 ;
  RECT 263.900 0.000 267.440 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 237.240 0.000 240.780 1.120 ;
  LAYER ME3 ;
  RECT 237.240 0.000 240.780 1.120 ;
  LAYER ME2 ;
  RECT 237.240 0.000 240.780 1.120 ;
  LAYER ME1 ;
  RECT 237.240 0.000 240.780 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 220.500 0.000 224.040 1.120 ;
  LAYER ME3 ;
  RECT 220.500 0.000 224.040 1.120 ;
  LAYER ME2 ;
  RECT 220.500 0.000 224.040 1.120 ;
  LAYER ME1 ;
  RECT 220.500 0.000 224.040 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 121.920 0.000 125.460 1.120 ;
  LAYER ME3 ;
  RECT 121.920 0.000 125.460 1.120 ;
  LAYER ME2 ;
  RECT 121.920 0.000 125.460 1.120 ;
  LAYER ME1 ;
  RECT 121.920 0.000 125.460 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 100.220 0.000 103.760 1.120 ;
  LAYER ME3 ;
  RECT 100.220 0.000 103.760 1.120 ;
  LAYER ME2 ;
  RECT 100.220 0.000 103.760 1.120 ;
  LAYER ME1 ;
  RECT 100.220 0.000 103.760 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 83.480 0.000 87.020 1.120 ;
  LAYER ME3 ;
  RECT 83.480 0.000 87.020 1.120 ;
  LAYER ME2 ;
  RECT 83.480 0.000 87.020 1.120 ;
  LAYER ME1 ;
  RECT 83.480 0.000 87.020 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 56.820 0.000 60.360 1.120 ;
  LAYER ME3 ;
  RECT 56.820 0.000 60.360 1.120 ;
  LAYER ME2 ;
  RECT 56.820 0.000 60.360 1.120 ;
  LAYER ME1 ;
  RECT 56.820 0.000 60.360 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER ME3 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER ME2 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER ME1 ;
  RECT 35.740 0.000 39.280 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER ME3 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER ME2 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER ME1 ;
  RECT 14.040 0.000 17.580 1.120 ;
 END
END VCC
PIN GND
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
 PORT
  LAYER ME4 ;
  RECT 325.620 278.660 326.740 281.900 ;
  LAYER ME3 ;
  RECT 325.620 278.660 326.740 281.900 ;
  LAYER ME2 ;
  RECT 325.620 278.660 326.740 281.900 ;
  LAYER ME1 ;
  RECT 325.620 278.660 326.740 281.900 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.620 270.820 326.740 274.060 ;
  LAYER ME3 ;
  RECT 325.620 270.820 326.740 274.060 ;
  LAYER ME2 ;
  RECT 325.620 270.820 326.740 274.060 ;
  LAYER ME1 ;
  RECT 325.620 270.820 326.740 274.060 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.620 262.980 326.740 266.220 ;
  LAYER ME3 ;
  RECT 325.620 262.980 326.740 266.220 ;
  LAYER ME2 ;
  RECT 325.620 262.980 326.740 266.220 ;
  LAYER ME1 ;
  RECT 325.620 262.980 326.740 266.220 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.620 255.140 326.740 258.380 ;
  LAYER ME3 ;
  RECT 325.620 255.140 326.740 258.380 ;
  LAYER ME2 ;
  RECT 325.620 255.140 326.740 258.380 ;
  LAYER ME1 ;
  RECT 325.620 255.140 326.740 258.380 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.620 247.300 326.740 250.540 ;
  LAYER ME3 ;
  RECT 325.620 247.300 326.740 250.540 ;
  LAYER ME2 ;
  RECT 325.620 247.300 326.740 250.540 ;
  LAYER ME1 ;
  RECT 325.620 247.300 326.740 250.540 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.620 208.100 326.740 211.340 ;
  LAYER ME3 ;
  RECT 325.620 208.100 326.740 211.340 ;
  LAYER ME2 ;
  RECT 325.620 208.100 326.740 211.340 ;
  LAYER ME1 ;
  RECT 325.620 208.100 326.740 211.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.620 200.260 326.740 203.500 ;
  LAYER ME3 ;
  RECT 325.620 200.260 326.740 203.500 ;
  LAYER ME2 ;
  RECT 325.620 200.260 326.740 203.500 ;
  LAYER ME1 ;
  RECT 325.620 200.260 326.740 203.500 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.620 192.420 326.740 195.660 ;
  LAYER ME3 ;
  RECT 325.620 192.420 326.740 195.660 ;
  LAYER ME2 ;
  RECT 325.620 192.420 326.740 195.660 ;
  LAYER ME1 ;
  RECT 325.620 192.420 326.740 195.660 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.620 184.580 326.740 187.820 ;
  LAYER ME3 ;
  RECT 325.620 184.580 326.740 187.820 ;
  LAYER ME2 ;
  RECT 325.620 184.580 326.740 187.820 ;
  LAYER ME1 ;
  RECT 325.620 184.580 326.740 187.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.620 176.740 326.740 179.980 ;
  LAYER ME3 ;
  RECT 325.620 176.740 326.740 179.980 ;
  LAYER ME2 ;
  RECT 325.620 176.740 326.740 179.980 ;
  LAYER ME1 ;
  RECT 325.620 176.740 326.740 179.980 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.620 168.900 326.740 172.140 ;
  LAYER ME3 ;
  RECT 325.620 168.900 326.740 172.140 ;
  LAYER ME2 ;
  RECT 325.620 168.900 326.740 172.140 ;
  LAYER ME1 ;
  RECT 325.620 168.900 326.740 172.140 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.620 129.700 326.740 132.940 ;
  LAYER ME3 ;
  RECT 325.620 129.700 326.740 132.940 ;
  LAYER ME2 ;
  RECT 325.620 129.700 326.740 132.940 ;
  LAYER ME1 ;
  RECT 325.620 129.700 326.740 132.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.620 121.860 326.740 125.100 ;
  LAYER ME3 ;
  RECT 325.620 121.860 326.740 125.100 ;
  LAYER ME2 ;
  RECT 325.620 121.860 326.740 125.100 ;
  LAYER ME1 ;
  RECT 325.620 121.860 326.740 125.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.620 114.020 326.740 117.260 ;
  LAYER ME3 ;
  RECT 325.620 114.020 326.740 117.260 ;
  LAYER ME2 ;
  RECT 325.620 114.020 326.740 117.260 ;
  LAYER ME1 ;
  RECT 325.620 114.020 326.740 117.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.620 106.180 326.740 109.420 ;
  LAYER ME3 ;
  RECT 325.620 106.180 326.740 109.420 ;
  LAYER ME2 ;
  RECT 325.620 106.180 326.740 109.420 ;
  LAYER ME1 ;
  RECT 325.620 106.180 326.740 109.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.620 98.340 326.740 101.580 ;
  LAYER ME3 ;
  RECT 325.620 98.340 326.740 101.580 ;
  LAYER ME2 ;
  RECT 325.620 98.340 326.740 101.580 ;
  LAYER ME1 ;
  RECT 325.620 98.340 326.740 101.580 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.620 90.500 326.740 93.740 ;
  LAYER ME3 ;
  RECT 325.620 90.500 326.740 93.740 ;
  LAYER ME2 ;
  RECT 325.620 90.500 326.740 93.740 ;
  LAYER ME1 ;
  RECT 325.620 90.500 326.740 93.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.620 51.300 326.740 54.540 ;
  LAYER ME3 ;
  RECT 325.620 51.300 326.740 54.540 ;
  LAYER ME2 ;
  RECT 325.620 51.300 326.740 54.540 ;
  LAYER ME1 ;
  RECT 325.620 51.300 326.740 54.540 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.620 43.460 326.740 46.700 ;
  LAYER ME3 ;
  RECT 325.620 43.460 326.740 46.700 ;
  LAYER ME2 ;
  RECT 325.620 43.460 326.740 46.700 ;
  LAYER ME1 ;
  RECT 325.620 43.460 326.740 46.700 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.620 35.620 326.740 38.860 ;
  LAYER ME3 ;
  RECT 325.620 35.620 326.740 38.860 ;
  LAYER ME2 ;
  RECT 325.620 35.620 326.740 38.860 ;
  LAYER ME1 ;
  RECT 325.620 35.620 326.740 38.860 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.620 27.780 326.740 31.020 ;
  LAYER ME3 ;
  RECT 325.620 27.780 326.740 31.020 ;
  LAYER ME2 ;
  RECT 325.620 27.780 326.740 31.020 ;
  LAYER ME1 ;
  RECT 325.620 27.780 326.740 31.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.620 19.940 326.740 23.180 ;
  LAYER ME3 ;
  RECT 325.620 19.940 326.740 23.180 ;
  LAYER ME2 ;
  RECT 325.620 19.940 326.740 23.180 ;
  LAYER ME1 ;
  RECT 325.620 19.940 326.740 23.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.620 12.100 326.740 15.340 ;
  LAYER ME3 ;
  RECT 325.620 12.100 326.740 15.340 ;
  LAYER ME2 ;
  RECT 325.620 12.100 326.740 15.340 ;
  LAYER ME1 ;
  RECT 325.620 12.100 326.740 15.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 278.660 1.120 281.900 ;
  LAYER ME3 ;
  RECT 0.000 278.660 1.120 281.900 ;
  LAYER ME2 ;
  RECT 0.000 278.660 1.120 281.900 ;
  LAYER ME1 ;
  RECT 0.000 278.660 1.120 281.900 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 270.820 1.120 274.060 ;
  LAYER ME3 ;
  RECT 0.000 270.820 1.120 274.060 ;
  LAYER ME2 ;
  RECT 0.000 270.820 1.120 274.060 ;
  LAYER ME1 ;
  RECT 0.000 270.820 1.120 274.060 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 262.980 1.120 266.220 ;
  LAYER ME3 ;
  RECT 0.000 262.980 1.120 266.220 ;
  LAYER ME2 ;
  RECT 0.000 262.980 1.120 266.220 ;
  LAYER ME1 ;
  RECT 0.000 262.980 1.120 266.220 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 255.140 1.120 258.380 ;
  LAYER ME3 ;
  RECT 0.000 255.140 1.120 258.380 ;
  LAYER ME2 ;
  RECT 0.000 255.140 1.120 258.380 ;
  LAYER ME1 ;
  RECT 0.000 255.140 1.120 258.380 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 247.300 1.120 250.540 ;
  LAYER ME3 ;
  RECT 0.000 247.300 1.120 250.540 ;
  LAYER ME2 ;
  RECT 0.000 247.300 1.120 250.540 ;
  LAYER ME1 ;
  RECT 0.000 247.300 1.120 250.540 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 208.100 1.120 211.340 ;
  LAYER ME3 ;
  RECT 0.000 208.100 1.120 211.340 ;
  LAYER ME2 ;
  RECT 0.000 208.100 1.120 211.340 ;
  LAYER ME1 ;
  RECT 0.000 208.100 1.120 211.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 200.260 1.120 203.500 ;
  LAYER ME3 ;
  RECT 0.000 200.260 1.120 203.500 ;
  LAYER ME2 ;
  RECT 0.000 200.260 1.120 203.500 ;
  LAYER ME1 ;
  RECT 0.000 200.260 1.120 203.500 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 192.420 1.120 195.660 ;
  LAYER ME3 ;
  RECT 0.000 192.420 1.120 195.660 ;
  LAYER ME2 ;
  RECT 0.000 192.420 1.120 195.660 ;
  LAYER ME1 ;
  RECT 0.000 192.420 1.120 195.660 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 184.580 1.120 187.820 ;
  LAYER ME3 ;
  RECT 0.000 184.580 1.120 187.820 ;
  LAYER ME2 ;
  RECT 0.000 184.580 1.120 187.820 ;
  LAYER ME1 ;
  RECT 0.000 184.580 1.120 187.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 176.740 1.120 179.980 ;
  LAYER ME3 ;
  RECT 0.000 176.740 1.120 179.980 ;
  LAYER ME2 ;
  RECT 0.000 176.740 1.120 179.980 ;
  LAYER ME1 ;
  RECT 0.000 176.740 1.120 179.980 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 168.900 1.120 172.140 ;
  LAYER ME3 ;
  RECT 0.000 168.900 1.120 172.140 ;
  LAYER ME2 ;
  RECT 0.000 168.900 1.120 172.140 ;
  LAYER ME1 ;
  RECT 0.000 168.900 1.120 172.140 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER ME3 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER ME2 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER ME1 ;
  RECT 0.000 129.700 1.120 132.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER ME3 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER ME2 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER ME1 ;
  RECT 0.000 121.860 1.120 125.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER ME3 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER ME2 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER ME1 ;
  RECT 0.000 114.020 1.120 117.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER ME3 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER ME2 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER ME1 ;
  RECT 0.000 106.180 1.120 109.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER ME3 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER ME2 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER ME1 ;
  RECT 0.000 98.340 1.120 101.580 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER ME3 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER ME2 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER ME1 ;
  RECT 0.000 90.500 1.120 93.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER ME3 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER ME2 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER ME1 ;
  RECT 0.000 51.300 1.120 54.540 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER ME3 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER ME2 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER ME1 ;
  RECT 0.000 43.460 1.120 46.700 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER ME3 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER ME2 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER ME1 ;
  RECT 0.000 35.620 1.120 38.860 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER ME3 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER ME2 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER ME1 ;
  RECT 0.000 27.780 1.120 31.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER ME3 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER ME2 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER ME1 ;
  RECT 0.000 19.940 1.120 23.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER ME3 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER ME2 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER ME1 ;
  RECT 0.000 12.100 1.120 15.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 307.300 292.880 310.840 294.000 ;
  LAYER ME3 ;
  RECT 307.300 292.880 310.840 294.000 ;
  LAYER ME2 ;
  RECT 307.300 292.880 310.840 294.000 ;
  LAYER ME1 ;
  RECT 307.300 292.880 310.840 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 298.620 292.880 302.160 294.000 ;
  LAYER ME3 ;
  RECT 298.620 292.880 302.160 294.000 ;
  LAYER ME2 ;
  RECT 298.620 292.880 302.160 294.000 ;
  LAYER ME1 ;
  RECT 298.620 292.880 302.160 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 289.940 292.880 293.480 294.000 ;
  LAYER ME3 ;
  RECT 289.940 292.880 293.480 294.000 ;
  LAYER ME2 ;
  RECT 289.940 292.880 293.480 294.000 ;
  LAYER ME1 ;
  RECT 289.940 292.880 293.480 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 281.260 292.880 284.800 294.000 ;
  LAYER ME3 ;
  RECT 281.260 292.880 284.800 294.000 ;
  LAYER ME2 ;
  RECT 281.260 292.880 284.800 294.000 ;
  LAYER ME1 ;
  RECT 281.260 292.880 284.800 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 272.580 292.880 276.120 294.000 ;
  LAYER ME3 ;
  RECT 272.580 292.880 276.120 294.000 ;
  LAYER ME2 ;
  RECT 272.580 292.880 276.120 294.000 ;
  LAYER ME1 ;
  RECT 272.580 292.880 276.120 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 229.180 292.880 232.720 294.000 ;
  LAYER ME3 ;
  RECT 229.180 292.880 232.720 294.000 ;
  LAYER ME2 ;
  RECT 229.180 292.880 232.720 294.000 ;
  LAYER ME1 ;
  RECT 229.180 292.880 232.720 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 220.500 292.880 224.040 294.000 ;
  LAYER ME3 ;
  RECT 220.500 292.880 224.040 294.000 ;
  LAYER ME2 ;
  RECT 220.500 292.880 224.040 294.000 ;
  LAYER ME1 ;
  RECT 220.500 292.880 224.040 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 211.820 292.880 215.360 294.000 ;
  LAYER ME3 ;
  RECT 211.820 292.880 215.360 294.000 ;
  LAYER ME2 ;
  RECT 211.820 292.880 215.360 294.000 ;
  LAYER ME1 ;
  RECT 211.820 292.880 215.360 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 203.140 292.880 206.680 294.000 ;
  LAYER ME3 ;
  RECT 203.140 292.880 206.680 294.000 ;
  LAYER ME2 ;
  RECT 203.140 292.880 206.680 294.000 ;
  LAYER ME1 ;
  RECT 203.140 292.880 206.680 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 194.460 292.880 198.000 294.000 ;
  LAYER ME3 ;
  RECT 194.460 292.880 198.000 294.000 ;
  LAYER ME2 ;
  RECT 194.460 292.880 198.000 294.000 ;
  LAYER ME1 ;
  RECT 194.460 292.880 198.000 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 185.780 292.880 189.320 294.000 ;
  LAYER ME3 ;
  RECT 185.780 292.880 189.320 294.000 ;
  LAYER ME2 ;
  RECT 185.780 292.880 189.320 294.000 ;
  LAYER ME1 ;
  RECT 185.780 292.880 189.320 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 142.380 292.880 145.920 294.000 ;
  LAYER ME3 ;
  RECT 142.380 292.880 145.920 294.000 ;
  LAYER ME2 ;
  RECT 142.380 292.880 145.920 294.000 ;
  LAYER ME1 ;
  RECT 142.380 292.880 145.920 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 133.700 292.880 137.240 294.000 ;
  LAYER ME3 ;
  RECT 133.700 292.880 137.240 294.000 ;
  LAYER ME2 ;
  RECT 133.700 292.880 137.240 294.000 ;
  LAYER ME1 ;
  RECT 133.700 292.880 137.240 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 125.020 292.880 128.560 294.000 ;
  LAYER ME3 ;
  RECT 125.020 292.880 128.560 294.000 ;
  LAYER ME2 ;
  RECT 125.020 292.880 128.560 294.000 ;
  LAYER ME1 ;
  RECT 125.020 292.880 128.560 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 116.340 292.880 119.880 294.000 ;
  LAYER ME3 ;
  RECT 116.340 292.880 119.880 294.000 ;
  LAYER ME2 ;
  RECT 116.340 292.880 119.880 294.000 ;
  LAYER ME1 ;
  RECT 116.340 292.880 119.880 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 107.660 292.880 111.200 294.000 ;
  LAYER ME3 ;
  RECT 107.660 292.880 111.200 294.000 ;
  LAYER ME2 ;
  RECT 107.660 292.880 111.200 294.000 ;
  LAYER ME1 ;
  RECT 107.660 292.880 111.200 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 98.980 292.880 102.520 294.000 ;
  LAYER ME3 ;
  RECT 98.980 292.880 102.520 294.000 ;
  LAYER ME2 ;
  RECT 98.980 292.880 102.520 294.000 ;
  LAYER ME1 ;
  RECT 98.980 292.880 102.520 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 55.580 292.880 59.120 294.000 ;
  LAYER ME3 ;
  RECT 55.580 292.880 59.120 294.000 ;
  LAYER ME2 ;
  RECT 55.580 292.880 59.120 294.000 ;
  LAYER ME1 ;
  RECT 55.580 292.880 59.120 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 46.900 292.880 50.440 294.000 ;
  LAYER ME3 ;
  RECT 46.900 292.880 50.440 294.000 ;
  LAYER ME2 ;
  RECT 46.900 292.880 50.440 294.000 ;
  LAYER ME1 ;
  RECT 46.900 292.880 50.440 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 38.220 292.880 41.760 294.000 ;
  LAYER ME3 ;
  RECT 38.220 292.880 41.760 294.000 ;
  LAYER ME2 ;
  RECT 38.220 292.880 41.760 294.000 ;
  LAYER ME1 ;
  RECT 38.220 292.880 41.760 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 29.540 292.880 33.080 294.000 ;
  LAYER ME3 ;
  RECT 29.540 292.880 33.080 294.000 ;
  LAYER ME2 ;
  RECT 29.540 292.880 33.080 294.000 ;
  LAYER ME1 ;
  RECT 29.540 292.880 33.080 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 20.860 292.880 24.400 294.000 ;
  LAYER ME3 ;
  RECT 20.860 292.880 24.400 294.000 ;
  LAYER ME2 ;
  RECT 20.860 292.880 24.400 294.000 ;
  LAYER ME1 ;
  RECT 20.860 292.880 24.400 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 12.180 292.880 15.720 294.000 ;
  LAYER ME3 ;
  RECT 12.180 292.880 15.720 294.000 ;
  LAYER ME2 ;
  RECT 12.180 292.880 15.720 294.000 ;
  LAYER ME1 ;
  RECT 12.180 292.880 15.720 294.000 ;
 END
 PORT
  LAYER ME4 ;
  RECT 315.360 0.000 318.900 1.120 ;
  LAYER ME3 ;
  RECT 315.360 0.000 318.900 1.120 ;
  LAYER ME2 ;
  RECT 315.360 0.000 318.900 1.120 ;
  LAYER ME1 ;
  RECT 315.360 0.000 318.900 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 293.660 0.000 297.200 1.120 ;
  LAYER ME3 ;
  RECT 293.660 0.000 297.200 1.120 ;
  LAYER ME2 ;
  RECT 293.660 0.000 297.200 1.120 ;
  LAYER ME1 ;
  RECT 293.660 0.000 297.200 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 276.920 0.000 280.460 1.120 ;
  LAYER ME3 ;
  RECT 276.920 0.000 280.460 1.120 ;
  LAYER ME2 ;
  RECT 276.920 0.000 280.460 1.120 ;
  LAYER ME1 ;
  RECT 276.920 0.000 280.460 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 250.880 0.000 254.420 1.120 ;
  LAYER ME3 ;
  RECT 250.880 0.000 254.420 1.120 ;
  LAYER ME2 ;
  RECT 250.880 0.000 254.420 1.120 ;
  LAYER ME1 ;
  RECT 250.880 0.000 254.420 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 229.180 0.000 232.720 1.120 ;
  LAYER ME3 ;
  RECT 229.180 0.000 232.720 1.120 ;
  LAYER ME2 ;
  RECT 229.180 0.000 232.720 1.120 ;
  LAYER ME1 ;
  RECT 229.180 0.000 232.720 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 126.260 0.000 129.800 1.120 ;
  LAYER ME3 ;
  RECT 126.260 0.000 129.800 1.120 ;
  LAYER ME2 ;
  RECT 126.260 0.000 129.800 1.120 ;
  LAYER ME1 ;
  RECT 126.260 0.000 129.800 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 113.860 0.000 117.400 1.120 ;
  LAYER ME3 ;
  RECT 113.860 0.000 117.400 1.120 ;
  LAYER ME2 ;
  RECT 113.860 0.000 117.400 1.120 ;
  LAYER ME1 ;
  RECT 113.860 0.000 117.400 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 92.160 0.000 95.700 1.120 ;
  LAYER ME3 ;
  RECT 92.160 0.000 95.700 1.120 ;
  LAYER ME2 ;
  RECT 92.160 0.000 95.700 1.120 ;
  LAYER ME1 ;
  RECT 92.160 0.000 95.700 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER ME3 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER ME2 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER ME1 ;
  RECT 70.460 0.000 74.000 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 43.800 0.000 47.340 1.120 ;
  LAYER ME3 ;
  RECT 43.800 0.000 47.340 1.120 ;
  LAYER ME2 ;
  RECT 43.800 0.000 47.340 1.120 ;
  LAYER ME1 ;
  RECT 43.800 0.000 47.340 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER ME3 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER ME2 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER ME1 ;
  RECT 27.060 0.000 30.600 1.120 ;
 END
END GND
PIN DO15
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 313.160 0.000 314.280 1.120 ;
  LAYER ME3 ;
  RECT 313.160 0.000 314.280 1.120 ;
  LAYER ME2 ;
  RECT 313.160 0.000 314.280 1.120 ;
  LAYER ME1 ;
  RECT 313.160 0.000 314.280 1.120 ;
 END
END DO15
PIN DI15
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 305.100 0.000 306.220 1.120 ;
  LAYER ME3 ;
  RECT 305.100 0.000 306.220 1.120 ;
  LAYER ME2 ;
  RECT 305.100 0.000 306.220 1.120 ;
  LAYER ME1 ;
  RECT 305.100 0.000 306.220 1.120 ;
 END
END DI15
PIN DO14
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 300.140 0.000 301.260 1.120 ;
  LAYER ME3 ;
  RECT 300.140 0.000 301.260 1.120 ;
  LAYER ME2 ;
  RECT 300.140 0.000 301.260 1.120 ;
  LAYER ME1 ;
  RECT 300.140 0.000 301.260 1.120 ;
 END
END DO14
PIN DI14
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 291.460 0.000 292.580 1.120 ;
  LAYER ME3 ;
  RECT 291.460 0.000 292.580 1.120 ;
  LAYER ME2 ;
  RECT 291.460 0.000 292.580 1.120 ;
  LAYER ME1 ;
  RECT 291.460 0.000 292.580 1.120 ;
 END
END DI14
PIN DO13
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 283.400 0.000 284.520 1.120 ;
  LAYER ME3 ;
  RECT 283.400 0.000 284.520 1.120 ;
  LAYER ME2 ;
  RECT 283.400 0.000 284.520 1.120 ;
  LAYER ME1 ;
  RECT 283.400 0.000 284.520 1.120 ;
 END
END DO13
PIN DI13
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 274.720 0.000 275.840 1.120 ;
  LAYER ME3 ;
  RECT 274.720 0.000 275.840 1.120 ;
  LAYER ME2 ;
  RECT 274.720 0.000 275.840 1.120 ;
  LAYER ME1 ;
  RECT 274.720 0.000 275.840 1.120 ;
 END
END DI13
PIN DO12
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 270.380 0.000 271.500 1.120 ;
  LAYER ME3 ;
  RECT 270.380 0.000 271.500 1.120 ;
  LAYER ME2 ;
  RECT 270.380 0.000 271.500 1.120 ;
  LAYER ME1 ;
  RECT 270.380 0.000 271.500 1.120 ;
 END
END DO12
PIN DI12
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 261.700 0.000 262.820 1.120 ;
  LAYER ME3 ;
  RECT 261.700 0.000 262.820 1.120 ;
  LAYER ME2 ;
  RECT 261.700 0.000 262.820 1.120 ;
  LAYER ME1 ;
  RECT 261.700 0.000 262.820 1.120 ;
 END
END DI12
PIN DO11
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 256.740 0.000 257.860 1.120 ;
  LAYER ME3 ;
  RECT 256.740 0.000 257.860 1.120 ;
  LAYER ME2 ;
  RECT 256.740 0.000 257.860 1.120 ;
  LAYER ME1 ;
  RECT 256.740 0.000 257.860 1.120 ;
 END
END DO11
PIN DI11
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 248.680 0.000 249.800 1.120 ;
  LAYER ME3 ;
  RECT 248.680 0.000 249.800 1.120 ;
  LAYER ME2 ;
  RECT 248.680 0.000 249.800 1.120 ;
  LAYER ME1 ;
  RECT 248.680 0.000 249.800 1.120 ;
 END
END DI11
PIN DO10
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 243.720 0.000 244.840 1.120 ;
  LAYER ME3 ;
  RECT 243.720 0.000 244.840 1.120 ;
  LAYER ME2 ;
  RECT 243.720 0.000 244.840 1.120 ;
  LAYER ME1 ;
  RECT 243.720 0.000 244.840 1.120 ;
 END
END DO10
PIN DI10
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 235.040 0.000 236.160 1.120 ;
  LAYER ME3 ;
  RECT 235.040 0.000 236.160 1.120 ;
  LAYER ME2 ;
  RECT 235.040 0.000 236.160 1.120 ;
  LAYER ME1 ;
  RECT 235.040 0.000 236.160 1.120 ;
 END
END DI10
PIN DO9
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 226.980 0.000 228.100 1.120 ;
  LAYER ME3 ;
  RECT 226.980 0.000 228.100 1.120 ;
  LAYER ME2 ;
  RECT 226.980 0.000 228.100 1.120 ;
  LAYER ME1 ;
  RECT 226.980 0.000 228.100 1.120 ;
 END
END DO9
PIN DI9
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 218.300 0.000 219.420 1.120 ;
  LAYER ME3 ;
  RECT 218.300 0.000 219.420 1.120 ;
  LAYER ME2 ;
  RECT 218.300 0.000 219.420 1.120 ;
  LAYER ME1 ;
  RECT 218.300 0.000 219.420 1.120 ;
 END
END DI9
PIN DO8
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 213.340 0.000 214.460 1.120 ;
  LAYER ME3 ;
  RECT 213.340 0.000 214.460 1.120 ;
  LAYER ME2 ;
  RECT 213.340 0.000 214.460 1.120 ;
  LAYER ME1 ;
  RECT 213.340 0.000 214.460 1.120 ;
 END
END DO8
PIN DI8
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 205.280 0.000 206.400 1.120 ;
  LAYER ME3 ;
  RECT 205.280 0.000 206.400 1.120 ;
  LAYER ME2 ;
  RECT 205.280 0.000 206.400 1.120 ;
  LAYER ME1 ;
  RECT 205.280 0.000 206.400 1.120 ;
 END
END DI8
PIN A1
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 199.700 0.000 200.820 1.120 ;
  LAYER ME3 ;
  RECT 199.700 0.000 200.820 1.120 ;
  LAYER ME2 ;
  RECT 199.700 0.000 200.820 1.120 ;
  LAYER ME1 ;
  RECT 199.700 0.000 200.820 1.120 ;
 END
END A1
PIN WEB
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER ME4 ;
  RECT 197.840 0.000 198.960 1.120 ;
  LAYER ME3 ;
  RECT 197.840 0.000 198.960 1.120 ;
  LAYER ME2 ;
  RECT 197.840 0.000 198.960 1.120 ;
  LAYER ME1 ;
  RECT 197.840 0.000 198.960 1.120 ;
 END
END WEB
PIN OE
  DIRECTION INPUT ;
  CAPACITANCE 0.033 ;
 PORT
  LAYER ME4 ;
  RECT 192.880 0.000 194.000 1.120 ;
  LAYER ME3 ;
  RECT 192.880 0.000 194.000 1.120 ;
  LAYER ME2 ;
  RECT 192.880 0.000 194.000 1.120 ;
  LAYER ME1 ;
  RECT 192.880 0.000 194.000 1.120 ;
 END
END OE
PIN CS
  DIRECTION INPUT ;
  CAPACITANCE 0.123 ;
 PORT
  LAYER ME4 ;
  RECT 191.020 0.000 192.140 1.120 ;
  LAYER ME3 ;
  RECT 191.020 0.000 192.140 1.120 ;
  LAYER ME2 ;
  RECT 191.020 0.000 192.140 1.120 ;
  LAYER ME1 ;
  RECT 191.020 0.000 192.140 1.120 ;
 END
END CS
PIN A2
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 169.320 0.000 170.440 1.120 ;
  LAYER ME3 ;
  RECT 169.320 0.000 170.440 1.120 ;
  LAYER ME2 ;
  RECT 169.320 0.000 170.440 1.120 ;
  LAYER ME1 ;
  RECT 169.320 0.000 170.440 1.120 ;
 END
END A2
PIN CK
  DIRECTION INPUT ;
  CAPACITANCE 0.063 ;
 PORT
  LAYER ME4 ;
  RECT 166.220 0.000 167.340 1.120 ;
  LAYER ME3 ;
  RECT 166.220 0.000 167.340 1.120 ;
  LAYER ME2 ;
  RECT 166.220 0.000 167.340 1.120 ;
  LAYER ME1 ;
  RECT 166.220 0.000 167.340 1.120 ;
 END
END CK
PIN A0
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 163.740 0.000 164.860 1.120 ;
  LAYER ME3 ;
  RECT 163.740 0.000 164.860 1.120 ;
  LAYER ME2 ;
  RECT 163.740 0.000 164.860 1.120 ;
  LAYER ME1 ;
  RECT 163.740 0.000 164.860 1.120 ;
 END
END A0
PIN A3
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 160.020 0.000 161.140 1.120 ;
  LAYER ME3 ;
  RECT 160.020 0.000 161.140 1.120 ;
  LAYER ME2 ;
  RECT 160.020 0.000 161.140 1.120 ;
  LAYER ME1 ;
  RECT 160.020 0.000 161.140 1.120 ;
 END
END A3
PIN A4
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 151.960 0.000 153.080 1.120 ;
  LAYER ME3 ;
  RECT 151.960 0.000 153.080 1.120 ;
  LAYER ME2 ;
  RECT 151.960 0.000 153.080 1.120 ;
  LAYER ME1 ;
  RECT 151.960 0.000 153.080 1.120 ;
 END
END A4
PIN A5
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 148.860 0.000 149.980 1.120 ;
  LAYER ME3 ;
  RECT 148.860 0.000 149.980 1.120 ;
  LAYER ME2 ;
  RECT 148.860 0.000 149.980 1.120 ;
  LAYER ME1 ;
  RECT 148.860 0.000 149.980 1.120 ;
 END
END A5
PIN A6
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 141.420 0.000 142.540 1.120 ;
  LAYER ME3 ;
  RECT 141.420 0.000 142.540 1.120 ;
  LAYER ME2 ;
  RECT 141.420 0.000 142.540 1.120 ;
  LAYER ME1 ;
  RECT 141.420 0.000 142.540 1.120 ;
 END
END A6
PIN A7
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 138.320 0.000 139.440 1.120 ;
  LAYER ME3 ;
  RECT 138.320 0.000 139.440 1.120 ;
  LAYER ME2 ;
  RECT 138.320 0.000 139.440 1.120 ;
  LAYER ME1 ;
  RECT 138.320 0.000 139.440 1.120 ;
 END
END A7
PIN A8
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 130.880 0.000 132.000 1.120 ;
  LAYER ME3 ;
  RECT 130.880 0.000 132.000 1.120 ;
  LAYER ME2 ;
  RECT 130.880 0.000 132.000 1.120 ;
  LAYER ME1 ;
  RECT 130.880 0.000 132.000 1.120 ;
 END
END A8
PIN DO7
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 119.720 0.000 120.840 1.120 ;
  LAYER ME3 ;
  RECT 119.720 0.000 120.840 1.120 ;
  LAYER ME2 ;
  RECT 119.720 0.000 120.840 1.120 ;
  LAYER ME1 ;
  RECT 119.720 0.000 120.840 1.120 ;
 END
END DO7
PIN DI7
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 111.660 0.000 112.780 1.120 ;
  LAYER ME3 ;
  RECT 111.660 0.000 112.780 1.120 ;
  LAYER ME2 ;
  RECT 111.660 0.000 112.780 1.120 ;
  LAYER ME1 ;
  RECT 111.660 0.000 112.780 1.120 ;
 END
END DI7
PIN DO6
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER ME3 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER ME2 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER ME1 ;
  RECT 106.700 0.000 107.820 1.120 ;
 END
END DO6
PIN DI6
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 98.020 0.000 99.140 1.120 ;
  LAYER ME3 ;
  RECT 98.020 0.000 99.140 1.120 ;
  LAYER ME2 ;
  RECT 98.020 0.000 99.140 1.120 ;
  LAYER ME1 ;
  RECT 98.020 0.000 99.140 1.120 ;
 END
END DI6
PIN DO5
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 89.960 0.000 91.080 1.120 ;
  LAYER ME3 ;
  RECT 89.960 0.000 91.080 1.120 ;
  LAYER ME2 ;
  RECT 89.960 0.000 91.080 1.120 ;
  LAYER ME1 ;
  RECT 89.960 0.000 91.080 1.120 ;
 END
END DO5
PIN DI5
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 81.280 0.000 82.400 1.120 ;
  LAYER ME3 ;
  RECT 81.280 0.000 82.400 1.120 ;
  LAYER ME2 ;
  RECT 81.280 0.000 82.400 1.120 ;
  LAYER ME1 ;
  RECT 81.280 0.000 82.400 1.120 ;
 END
END DI5
PIN DO4
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 76.320 0.000 77.440 1.120 ;
  LAYER ME3 ;
  RECT 76.320 0.000 77.440 1.120 ;
  LAYER ME2 ;
  RECT 76.320 0.000 77.440 1.120 ;
  LAYER ME1 ;
  RECT 76.320 0.000 77.440 1.120 ;
 END
END DO4
PIN DI4
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 68.260 0.000 69.380 1.120 ;
  LAYER ME3 ;
  RECT 68.260 0.000 69.380 1.120 ;
  LAYER ME2 ;
  RECT 68.260 0.000 69.380 1.120 ;
  LAYER ME1 ;
  RECT 68.260 0.000 69.380 1.120 ;
 END
END DI4
PIN DO3
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 63.300 0.000 64.420 1.120 ;
  LAYER ME3 ;
  RECT 63.300 0.000 64.420 1.120 ;
  LAYER ME2 ;
  RECT 63.300 0.000 64.420 1.120 ;
  LAYER ME1 ;
  RECT 63.300 0.000 64.420 1.120 ;
 END
END DO3
PIN DI3
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 54.620 0.000 55.740 1.120 ;
  LAYER ME3 ;
  RECT 54.620 0.000 55.740 1.120 ;
  LAYER ME2 ;
  RECT 54.620 0.000 55.740 1.120 ;
  LAYER ME1 ;
  RECT 54.620 0.000 55.740 1.120 ;
 END
END DI3
PIN DO2
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 50.280 0.000 51.400 1.120 ;
  LAYER ME3 ;
  RECT 50.280 0.000 51.400 1.120 ;
  LAYER ME2 ;
  RECT 50.280 0.000 51.400 1.120 ;
  LAYER ME1 ;
  RECT 50.280 0.000 51.400 1.120 ;
 END
END DO2
PIN DI2
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 41.600 0.000 42.720 1.120 ;
  LAYER ME3 ;
  RECT 41.600 0.000 42.720 1.120 ;
  LAYER ME2 ;
  RECT 41.600 0.000 42.720 1.120 ;
  LAYER ME1 ;
  RECT 41.600 0.000 42.720 1.120 ;
 END
END DI2
PIN DO1
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER ME3 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER ME2 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER ME1 ;
  RECT 33.540 0.000 34.660 1.120 ;
 END
END DO1
PIN DI1
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER ME3 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER ME2 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER ME1 ;
  RECT 24.860 0.000 25.980 1.120 ;
 END
END DI1
PIN DO0
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER ME3 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER ME2 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER ME1 ;
  RECT 19.900 0.000 21.020 1.120 ;
 END
END DO0
PIN DI0
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER ME3 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER ME2 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER ME1 ;
  RECT 11.840 0.000 12.960 1.120 ;
 END
END DI0
OBS
  LAYER ME1 SPACING 0.280 ;
  RECT 0.000 0.140 326.740 294.000 ;
  LAYER ME2 SPACING 0.320 ;
  RECT 0.000 0.140 326.740 294.000 ;
  LAYER ME3 SPACING 0.320 ;
  RECT 0.000 0.140 326.740 294.000 ;
  LAYER ME4 SPACING 0.600 ;
  RECT 0.000 0.140 326.740 294.000 ;
  LAYER VI1 ;
  RECT 0.000 0.140 326.740 294.000 ;
  LAYER VI2 ;
  RECT 0.000 0.140 326.740 294.000 ;
  LAYER VI3 ;
  RECT 0.000 0.140 326.740 294.000 ;
END
END MEM1_1
END LIBRARY



